module lsp

// method: ‘textDocument/declaration’
// response: Location | []Location | []LocationLink | none
// request: TextDocumentPositionParams